Circuit RLC
V1 1 0 PULSE(0 1 0 0 0 10M 20M)
R1 1 2 10K
C1 2 0 100N
L1 2 3 10M
R 3 4 10
VIL 4 0 DC 0
.CONTROL
IC V(2)=0
TRAN 1U 20M
PRINT V(2) > export-5.txt
.ENDC
.END