Circuit RLC
V1 1 0 AC 1
R1 1 2 10K
C1 2 0 100N
L1 2 3 10M
R 3 0 10
.CONTROL
AC DEC 100 100 100K
PRINT VDB(2) VP(2) > export-3.txt
.ENDC
.END
