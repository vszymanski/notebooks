Circuit RLC
V1 1 0 AC 1
R1 1 2 10K
C1 2 0 100N
L1 2 3 10M
R 3 4 10
VIL 4 0 DC 0
.CONTROL
AC DEC 100 100 100K
PRINT I(VIL) > export-4.txt
.ENDC
.END
